`timescale 1ns/100ps

module tb_rca_36b;

	reg [35:0] 	A;
	reg [35:0] 	B;
	reg 			Cin;

	wire [35:0] S;
	wire 			Cout;
	
	rca_36b uud(S, Cout, A, B, Cin);
	
	initial begin		
		// Initialize A, B, Cin
		A		= 36'b000000000000000000000000000000000000;
		B		= 36'b000000000000000000000000000000000000;
		Cin	= 36'b000000000000000000000000000000000000;
		
		
		#10;
		A		= 36'b111111111111111111111111111111111111;
		B		= 36'b000000000000000000000000000000000000;
		Cin	= 36'b000000000000000000000000000000000001;
		
		#10;
		A		= 36'b111111111111111111111111111111111111;
		B		= 36'b000000000000000000000000000000000001;
		Cin	= 36'b000000000000000000000000000000000000;
		
		#10;
		A		= 36'b000000000000000000000000000000000011;
		B		= 36'b000000000000000000000000000000000001;
		Cin	= 36'b000000000000000000000000000000000001;
		
		#10;
		A		= 36'b000000000000000000000000000000000000;
		B		= 36'b111111111111111111111111111111111101;
		Cin	= 36'b000000000000000000000000000000000001;
		
		#10;
		A		= 36'b000000000000000000000000000000000001;
		B		= 36'b000000000000000000000000000000000010;
		Cin	= 36'b000000000000000000000000000000000001;
		
		#10;
		end
endmodule
